interface accum_if(input clk,
            input rst);
    logic [7:0] data;
	logic valid;
endinterface

