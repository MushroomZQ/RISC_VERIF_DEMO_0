`include "../verif/register_uvm_env/register_pkg.sv"

package testcase_pkg;
    import uvm_pkg::*;
    import register_uvm_env_pkg::*;

    `include "register_testcase.sv"
endpackage: testcase_pkg
